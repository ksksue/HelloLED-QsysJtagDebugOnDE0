// qsys_led.v

// Generated using ACDS version 11.1 173 at 2011.12.10.02:41:08

`timescale 1 ps / 1 ps
module qsys_led (
		output wire [31:0] led_export, // led.export
		input  wire        clk_clk     // clk.clk
	);

	wire         master_0_master_reset_reset;                                        // master_0:master_reset_reset -> [rst_controller:reset_in0, rst_controller:reset_in1]
	wire         master_0_master_waitrequest;                                        // master_0_master_translator:av_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_writedata;                                          // master_0:master_writedata -> master_0_master_translator:av_writedata
	wire  [31:0] master_0_master_address;                                            // master_0:master_address -> master_0_master_translator:av_address
	wire         master_0_master_write;                                              // master_0:master_write -> master_0_master_translator:av_write
	wire         master_0_master_read;                                               // master_0:master_read -> master_0_master_translator:av_read
	wire  [31:0] master_0_master_readdata;                                           // master_0_master_translator:av_readdata -> master_0:master_readdata
	wire   [3:0] master_0_master_byteenable;                                         // master_0:master_byteenable -> master_0_master_translator:av_byteenable
	wire         master_0_master_readdatavalid;                                      // master_0_master_translator:av_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_translator_avalon_universal_master_0_waitrequest;   // led_s1_translator:uav_waitrequest -> master_0_master_translator:uav_waitrequest
	wire   [2:0] master_0_master_translator_avalon_universal_master_0_burstcount;    // master_0_master_translator:uav_burstcount -> led_s1_translator:uav_burstcount
	wire  [31:0] master_0_master_translator_avalon_universal_master_0_writedata;     // master_0_master_translator:uav_writedata -> led_s1_translator:uav_writedata
	wire  [31:0] master_0_master_translator_avalon_universal_master_0_address;       // master_0_master_translator:uav_address -> led_s1_translator:uav_address
	wire         master_0_master_translator_avalon_universal_master_0_lock;          // master_0_master_translator:uav_lock -> led_s1_translator:uav_lock
	wire         master_0_master_translator_avalon_universal_master_0_write;         // master_0_master_translator:uav_write -> led_s1_translator:uav_write
	wire         master_0_master_translator_avalon_universal_master_0_read;          // master_0_master_translator:uav_read -> led_s1_translator:uav_read
	wire  [31:0] master_0_master_translator_avalon_universal_master_0_readdata;      // led_s1_translator:uav_readdata -> master_0_master_translator:uav_readdata
	wire         master_0_master_translator_avalon_universal_master_0_debugaccess;   // master_0_master_translator:uav_debugaccess -> led_s1_translator:uav_debugaccess
	wire   [3:0] master_0_master_translator_avalon_universal_master_0_byteenable;    // master_0_master_translator:uav_byteenable -> led_s1_translator:uav_byteenable
	wire         master_0_master_translator_avalon_universal_master_0_readdatavalid; // led_s1_translator:uav_readdatavalid -> master_0_master_translator:uav_readdatavalid
	wire  [31:0] led_s1_translator_avalon_anti_slave_0_writedata;                    // led_s1_translator:av_writedata -> led:writedata
	wire   [1:0] led_s1_translator_avalon_anti_slave_0_address;                      // led_s1_translator:av_address -> led:address
	wire         led_s1_translator_avalon_anti_slave_0_chipselect;                   // led_s1_translator:av_chipselect -> led:chipselect
	wire         led_s1_translator_avalon_anti_slave_0_write;                        // led_s1_translator:av_write -> led:write_n
	wire  [31:0] led_s1_translator_avalon_anti_slave_0_readdata;                     // led:readdata -> led_s1_translator:av_readdata
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [led:reset_n, led_s1_translator:reset, master_0:clk_reset_reset, master_0_master_translator:reset]

	qsys_led_led led (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (led_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_export)                                        // external_connection.export
	);

	qsys_led_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                        //          clk.clk
		.clk_reset_reset      (rst_controller_reset_out_reset), //    clk_reset.reset
		.master_address       (master_0_master_address),        //       master.address
		.master_readdata      (master_0_master_readdata),       //             .readdata
		.master_read          (master_0_master_read),           //             .read
		.master_write         (master_0_master_write),          //             .write
		.master_writedata     (master_0_master_writedata),      //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),    //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid),  //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),     //             .byteenable
		.master_reset_reset   (master_0_master_reset_reset)     // master_reset.reset
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) master_0_master_translator (
		.clk                   (clk_clk),                                                            //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address           (master_0_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (master_0_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (master_0_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (master_0_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (master_0_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (master_0_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (master_0_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (master_0_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (master_0_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (master_0_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (master_0_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (master_0_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (master_0_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (master_0_master_byteenable),                                         //                          .byteenable
		.av_read               (master_0_master_read),                                               //                          .read
		.av_readdata           (master_0_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (master_0_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (master_0_master_write),                                              //                          .write
		.av_writedata          (master_0_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_s1_translator (
		.clk                   (clk_clk),                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (master_0_master_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (master_0_master_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read              (master_0_master_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write             (master_0_master_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest       (master_0_master_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (master_0_master_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (master_0_master_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata          (master_0_master_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata         (master_0_master_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock              (master_0_master_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess       (master_0_master_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address            (led_s1_translator_avalon_anti_slave_0_address),                      //      avalon_anti_slave_0.address
		.av_write              (led_s1_translator_avalon_anti_slave_0_write),                        //                         .write
		.av_readdata           (led_s1_translator_avalon_anti_slave_0_readdata),                     //                         .readdata
		.av_writedata          (led_s1_translator_avalon_anti_slave_0_writedata),                    //                         .writedata
		.av_chipselect         (led_s1_translator_avalon_anti_slave_0_chipselect),                   //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (master_0_master_reset_reset),    // reset_in0.reset
		.reset_in1  (master_0_master_reset_reset),    // reset_in1.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
